magic
tech sky130A
timestamp 1753449410
<< pwell >>
rect -223 -155 223 155
<< nmos >>
rect -125 -50 125 50
<< ndiff >>
rect -154 44 -125 50
rect -154 -44 -148 44
rect -131 -44 -125 44
rect -154 -50 -125 -44
rect 125 44 154 50
rect 125 -44 131 44
rect 148 -44 154 44
rect 125 -50 154 -44
<< ndiffc >>
rect -148 -44 -131 44
rect 131 -44 148 44
<< psubdiff >>
rect -205 120 -157 137
rect 157 120 205 137
rect -205 89 -188 120
rect 188 89 205 120
rect -205 -120 -188 -89
rect 188 -120 205 -89
rect -205 -137 -157 -120
rect 157 -137 205 -120
<< psubdiffcont >>
rect -157 120 157 137
rect -205 -89 -188 89
rect 188 -89 205 89
rect -157 -137 157 -120
<< poly >>
rect -125 86 125 94
rect -125 69 -117 86
rect 117 69 125 86
rect -125 50 125 69
rect -125 -69 125 -50
rect -125 -86 -117 -69
rect 117 -86 125 -69
rect -125 -94 125 -86
<< polycont >>
rect -117 69 117 86
rect -117 -86 117 -69
<< locali >>
rect -205 120 -157 137
rect 157 120 205 137
rect -205 89 -188 120
rect 188 89 205 120
rect -125 69 -117 86
rect 117 69 125 86
rect -148 44 -131 52
rect -148 -52 -131 -44
rect 131 44 148 52
rect 131 -52 148 -44
rect -125 -86 -117 -69
rect 117 -86 125 -69
rect -205 -120 -188 -89
rect 188 -120 205 -89
rect -205 -137 -157 -120
rect 157 -137 205 -120
<< viali >>
rect -117 69 117 86
rect -148 -44 -131 44
rect 131 -44 148 44
rect -117 -86 117 -69
<< metal1 >>
rect -123 86 123 89
rect -123 69 -117 86
rect 117 69 123 86
rect -123 66 123 69
rect -151 44 -128 50
rect -151 -44 -148 44
rect -131 -44 -128 44
rect -151 -50 -128 -44
rect 128 44 151 50
rect 128 -44 131 44
rect 148 -44 151 44
rect 128 -50 151 -44
rect -123 -69 123 -66
rect -123 -86 -117 -69
rect 117 -86 123 -69
rect -123 -89 123 -86
<< properties >>
string FIXED_BBOX -196 -128 196 128
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 2.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
