magic
tech sky130A
timestamp 1753449410
<< pwell >>
rect -223 -130 223 130
<< nmos >>
rect -125 -25 125 25
<< ndiff >>
rect -154 19 -125 25
rect -154 -19 -148 19
rect -131 -19 -125 19
rect -154 -25 -125 -19
rect 125 19 154 25
rect 125 -19 131 19
rect 148 -19 154 19
rect 125 -25 154 -19
<< ndiffc >>
rect -148 -19 -131 19
rect 131 -19 148 19
<< psubdiff >>
rect -205 95 -157 112
rect 157 95 205 112
rect -205 64 -188 95
rect 188 64 205 95
rect -205 -95 -188 -64
rect 188 -95 205 -64
rect -205 -112 -157 -95
rect 157 -112 205 -95
<< psubdiffcont >>
rect -157 95 157 112
rect -205 -64 -188 64
rect 188 -64 205 64
rect -157 -112 157 -95
<< poly >>
rect -125 61 125 69
rect -125 44 -117 61
rect 117 44 125 61
rect -125 25 125 44
rect -125 -44 125 -25
rect -125 -61 -117 -44
rect 117 -61 125 -44
rect -125 -69 125 -61
<< polycont >>
rect -117 44 117 61
rect -117 -61 117 -44
<< locali >>
rect -205 95 -157 112
rect 157 95 205 112
rect -205 64 -188 95
rect 188 64 205 95
rect -125 44 -117 61
rect 117 44 125 61
rect -148 19 -131 27
rect -148 -27 -131 -19
rect 131 19 148 27
rect 131 -27 148 -19
rect -125 -61 -117 -44
rect 117 -61 125 -44
rect -205 -95 -188 -64
rect 188 -95 205 -64
rect -205 -112 -157 -95
rect 157 -112 205 -95
<< viali >>
rect -117 44 117 61
rect -148 -19 -131 19
rect 131 -19 148 19
rect -117 -61 117 -44
<< metal1 >>
rect -123 61 123 64
rect -123 44 -117 61
rect 117 44 123 61
rect -123 41 123 44
rect -151 19 -128 25
rect -151 -19 -148 19
rect -131 -19 -128 19
rect -151 -25 -128 -19
rect 128 19 151 25
rect 128 -19 131 19
rect 148 -19 151 19
rect 128 -25 151 -19
rect -123 -44 123 -41
rect -123 -61 -117 -44
rect 117 -61 123 -44
rect -123 -64 123 -61
<< properties >>
string FIXED_BBOX -196 -103 196 103
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.5 l 2.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
