magic
tech sky130A
magscale 1 2
timestamp 1753449410
<< nwell >>
rect -446 -2219 446 2219
<< pmos >>
rect -250 -2000 250 2000
<< pdiff >>
rect -308 1988 -250 2000
rect -308 -1988 -296 1988
rect -262 -1988 -250 1988
rect -308 -2000 -250 -1988
rect 250 1988 308 2000
rect 250 -1988 262 1988
rect 296 -1988 308 1988
rect 250 -2000 308 -1988
<< pdiffc >>
rect -296 -1988 -262 1988
rect 262 -1988 296 1988
<< nsubdiff >>
rect -410 2149 -314 2183
rect 314 2149 410 2183
rect -410 2087 -376 2149
rect 376 2087 410 2149
rect -410 -2149 -376 -2087
rect 376 -2149 410 -2087
rect -410 -2183 -314 -2149
rect 314 -2183 410 -2149
<< nsubdiffcont >>
rect -314 2149 314 2183
rect -410 -2087 -376 2087
rect 376 -2087 410 2087
rect -314 -2183 314 -2149
<< poly >>
rect -250 2081 250 2097
rect -250 2047 -234 2081
rect 234 2047 250 2081
rect -250 2000 250 2047
rect -250 -2047 250 -2000
rect -250 -2081 -234 -2047
rect 234 -2081 250 -2047
rect -250 -2097 250 -2081
<< polycont >>
rect -234 2047 234 2081
rect -234 -2081 234 -2047
<< locali >>
rect -410 2149 -314 2183
rect 314 2149 410 2183
rect -410 2087 -376 2149
rect 376 2087 410 2149
rect -250 2047 -234 2081
rect 234 2047 250 2081
rect -296 1988 -262 2004
rect -296 -2004 -262 -1988
rect 262 1988 296 2004
rect 262 -2004 296 -1988
rect -250 -2081 -234 -2047
rect 234 -2081 250 -2047
rect -410 -2149 -376 -2087
rect 376 -2149 410 -2087
rect -410 -2183 -314 -2149
rect 314 -2183 410 -2149
<< viali >>
rect -234 2047 234 2081
rect -296 -1988 -262 1988
rect 262 -1988 296 1988
rect -234 -2081 234 -2047
<< metal1 >>
rect -246 2081 246 2087
rect -246 2047 -234 2081
rect 234 2047 246 2081
rect -246 2041 246 2047
rect -302 1988 -256 2000
rect -302 -1988 -296 1988
rect -262 -1988 -256 1988
rect -302 -2000 -256 -1988
rect 256 1988 302 2000
rect 256 -1988 262 1988
rect 296 -1988 302 1988
rect 256 -2000 302 -1988
rect -246 -2047 246 -2041
rect -246 -2081 -234 -2047
rect 234 -2081 246 -2047
rect -246 -2087 246 -2081
<< properties >>
string FIXED_BBOX -393 -2166 393 2166
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 20.0 l 2.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 class mosfet compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0 ad {int((nf+1)/2) * W/nf * 0.29} as {int((nf+2)/2) * W/nf * 0.29} pd {2*int((nf+1)/2) * (W/nf + 0.29)} ps {2*int((nf+2)/2) * (W/nf + 0.29)} nrd {0.29 / W} nrs {0.29 / W} sa 0 sb 0 sd 0 mult 1
<< end >>
