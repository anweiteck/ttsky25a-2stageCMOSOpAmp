magic
tech sky130A
magscale 1 2
timestamp 1753538542
<< locali >>
rect 9632 3216 11984 3240
rect 9632 3122 9680 3216
rect 11546 3122 11984 3216
rect 9632 2898 11984 3122
rect 9632 2876 11992 2898
rect 11422 2350 11992 2876
rect 9638 1532 9890 1952
rect 9638 1220 11986 1532
rect 9638 838 9890 1220
rect 11422 838 11986 1220
rect 9638 716 12772 838
rect 9638 604 9710 716
rect 12694 604 12772 716
rect 9638 556 12772 604
<< viali >>
rect 9680 3122 11546 3216
rect 9710 604 12694 716
<< metal1 >>
rect 11970 3750 12108 6518
rect 11970 3612 12016 3750
rect 12100 3612 12110 3750
rect 9378 3238 9578 3284
rect 9378 3216 11558 3238
rect 9378 3122 9680 3216
rect 11546 3122 11558 3216
rect 9378 3114 10480 3122
rect 10616 3114 11412 3122
rect 9378 3096 11412 3114
rect 9378 3084 9578 3096
rect 9796 2852 11264 3012
rect 9796 2810 10478 2852
rect 9798 2710 9962 2810
rect 9798 2538 10000 2710
rect 9798 1858 9922 2538
rect 10040 2446 10478 2810
rect 10514 2712 10610 2714
rect 10514 2704 10620 2712
rect 10514 2568 10526 2704
rect 10610 2568 10620 2704
rect 10514 2540 10620 2568
rect 10524 2538 10620 2540
rect 10660 2708 10764 2712
rect 10660 2698 10784 2708
rect 10660 2528 10682 2698
rect 10780 2528 10790 2698
rect 10660 2510 10782 2528
rect 10660 2504 10764 2510
rect 9798 1688 10004 1858
rect 9822 1686 10004 1688
rect 10114 1848 10364 1976
rect 10516 1848 10616 1856
rect 10114 1702 10164 1848
rect 10302 1702 10364 1848
rect 10114 1580 10364 1702
rect 10514 1700 10524 1848
rect 10606 1700 10616 1848
rect 10516 1684 10616 1700
rect 10652 1848 10764 2504
rect 10826 2448 11264 2852
rect 11388 3004 11412 3096
rect 11522 3004 11558 3122
rect 11970 3066 12108 3612
rect 11388 2712 11558 3004
rect 11310 2538 11558 2712
rect 11940 2540 12108 3066
rect 12146 3498 12580 6610
rect 12146 3330 12252 3498
rect 12480 3330 12580 3498
rect 10908 1860 11158 1974
rect 11940 1966 12082 2540
rect 12146 2448 12580 3330
rect 12630 3214 12866 6468
rect 12630 3004 12694 3214
rect 12830 3004 12866 3214
rect 12630 2582 12866 3004
rect 11940 1928 12102 1966
rect 11940 1908 12116 1928
rect 11940 1868 12024 1908
rect 10652 1696 10784 1848
rect 10908 1714 10974 1860
rect 11112 1714 11158 1860
rect 10908 1578 11158 1714
rect 11304 1688 11490 1860
rect 11414 1544 11490 1688
rect 10698 1528 11490 1544
rect 10698 1440 10706 1528
rect 10800 1440 11490 1528
rect 10698 1436 11490 1440
rect 9392 1270 10496 1272
rect 11214 1270 11860 1290
rect 9392 1200 11860 1270
rect 9392 1192 11252 1200
rect 9392 1138 10496 1192
rect 9386 1120 10496 1138
rect 10848 1154 11252 1192
rect 9386 1070 9972 1120
rect 9386 992 9998 1070
rect 9386 938 9972 992
rect 10046 910 10478 1120
rect 10704 1070 10804 1084
rect 10596 1068 10674 1070
rect 10522 994 10674 1068
rect 9410 752 9610 754
rect 10594 752 10674 994
rect 10704 992 10724 1070
rect 10784 992 10804 1070
rect 10704 978 10804 992
rect 10848 912 11254 1154
rect 11306 994 11462 1068
rect 11384 752 11462 994
rect 11574 948 11860 1200
rect 11966 1048 12024 1868
rect 12100 1048 12116 1908
rect 11966 1010 12116 1048
rect 11966 986 12102 1010
rect 12150 948 12566 2050
rect 12708 1964 12884 1966
rect 12628 986 12884 1964
rect 11572 906 12566 948
rect 11572 796 12562 906
rect 12152 792 12562 796
rect 12708 752 12884 986
rect 9410 716 12884 752
rect 9410 604 9710 716
rect 12694 604 12884 716
rect 9410 558 12884 604
rect 9410 556 9654 558
rect 9410 554 9610 556
rect 10120 452 10362 496
rect 10120 306 10168 452
rect 10308 306 10362 452
rect 10120 266 10362 306
rect 10916 454 11158 490
rect 10916 308 10958 454
rect 11098 308 11158 454
rect 10916 260 11158 308
rect 11874 458 12116 506
rect 11874 312 11920 458
rect 12060 312 12116 458
rect 11874 276 12116 312
<< via1 >>
rect 12016 3612 12100 3750
rect 10480 3122 10616 3216
rect 11412 3122 11522 3214
rect 10480 3114 10616 3122
rect 10526 2568 10610 2704
rect 10682 2528 10780 2698
rect 10164 1702 10302 1848
rect 10524 1700 10606 1848
rect 11412 3004 11522 3122
rect 12252 3330 12480 3498
rect 12694 3004 12830 3214
rect 10974 1714 11112 1860
rect 10706 1440 10800 1528
rect 10724 992 10784 1070
rect 12024 1048 12100 1908
rect 10168 306 10308 452
rect 10958 308 11098 454
rect 11920 312 12060 458
<< metal2 >>
rect 11600 3750 12112 3764
rect 11600 3738 12016 3750
rect 11600 3620 11638 3738
rect 11770 3620 12016 3738
rect 11600 3612 12016 3620
rect 12100 3612 12112 3750
rect 11600 3588 12112 3612
rect 10688 3498 12572 3528
rect 10678 3330 12252 3498
rect 12480 3330 12572 3498
rect 10678 3280 12572 3330
rect 10678 3250 10838 3280
rect 10530 3226 10618 3230
rect 10470 3216 10640 3226
rect 10470 3114 10480 3216
rect 10616 3114 10640 3216
rect 10470 2704 10640 3114
rect 10470 2568 10526 2704
rect 10610 2568 10640 2704
rect 10470 2556 10640 2568
rect 10678 3214 10836 3250
rect 10678 3022 10698 3214
rect 10810 3022 10836 3214
rect 10678 2698 10836 3022
rect 11390 3214 12870 3244
rect 11390 3004 11412 3214
rect 11522 3004 12694 3214
rect 12830 3004 12870 3214
rect 11390 2976 12870 3004
rect 10678 2528 10682 2698
rect 10780 2528 10836 2698
rect 10678 2520 10836 2528
rect 10682 2518 10780 2520
rect 10120 1848 10362 1978
rect 10916 1860 11158 1972
rect 10524 1856 10606 1858
rect 10120 1702 10164 1848
rect 10302 1702 10362 1848
rect 10120 452 10362 1702
rect 10516 1848 10698 1856
rect 10516 1700 10524 1848
rect 10606 1700 10698 1848
rect 10516 1684 10698 1700
rect 10622 1538 10698 1684
rect 10916 1714 10974 1860
rect 11112 1714 11158 1860
rect 10622 1528 10802 1538
rect 10622 1440 10706 1528
rect 10800 1440 10802 1528
rect 10622 1436 10802 1440
rect 10704 1282 10802 1436
rect 10706 1070 10802 1282
rect 10706 992 10724 1070
rect 10784 992 10802 1070
rect 10706 978 10802 992
rect 10120 306 10168 452
rect 10308 306 10362 452
rect 10120 266 10362 306
rect 10916 454 11158 1714
rect 10916 308 10958 454
rect 11098 308 11158 454
rect 10916 260 11158 308
rect 11876 1908 12118 1988
rect 11876 1048 12024 1908
rect 12100 1048 12118 1908
rect 11876 458 12118 1048
rect 11876 312 11920 458
rect 12060 312 12118 458
rect 11876 276 12118 312
<< via2 >>
rect 11638 3620 11770 3738
rect 10698 3022 10810 3214
<< metal3 >>
rect 7520 3780 11576 7556
rect 7520 3738 11838 3780
rect 7520 3620 11638 3738
rect 11770 3620 11838 3738
rect 7520 3546 11838 3620
rect 7520 3500 11576 3546
rect 10682 3214 10834 3222
rect 10682 3022 10698 3214
rect 10812 3022 10834 3214
rect 10682 3008 10834 3022
<< via3 >>
rect 10698 3022 10810 3214
rect 10810 3022 10812 3214
<< mimcap >>
rect 7548 3894 11548 7528
rect 7548 3660 10542 3894
rect 10780 3660 11548 3894
rect 7548 3528 11548 3660
<< mimcapcontact >>
rect 10542 3660 10780 3894
<< metal4 >>
rect 10506 3894 10804 3930
rect 10506 3660 10542 3894
rect 10780 3660 10804 3894
rect 10506 3500 10804 3660
rect 10686 3215 10804 3500
rect 10686 3214 10813 3215
rect 10686 3022 10698 3214
rect 10812 3022 10813 3214
rect 10686 3021 10813 3022
rect 10686 3016 10804 3021
use sky130_fd_pr__nfet_01v8_WH8SLP  XM1
timestamp 1753449410
transform 1 0 10264 0 1 1772
box -446 -310 446 310
use sky130_fd_pr__nfet_01v8_WH8SLP  XM2
timestamp 1753449410
transform 1 0 11050 0 1 1772
box -446 -310 446 310
use sky130_fd_pr__pfet_01v8_CQSGDB  XM3
timestamp 1753449410
transform 1 0 10262 0 1 2625
box -446 -319 446 319
use sky130_fd_pr__pfet_01v8_CQSGDB  XM4
timestamp 1753449410
transform 1 0 11048 0 1 2625
box -446 -319 446 319
use sky130_fd_pr__nfet_01v8_KW7QXQ  XM5
timestamp 1753449410
transform 1 0 11046 0 1 1032
box -446 -260 446 260
use sky130_fd_pr__pfet_01v8_AT44HV  XM6
timestamp 1753449410
transform 1 0 12368 0 1 4529
box -446 -2219 446 2219
use sky130_fd_pr__nfet_01v8_P9E9M2  XM7
timestamp 1753449410
transform 1 0 12364 0 1 1478
box -446 -710 446 710
use sky130_fd_pr__nfet_01v8_KW7QXQ  XM8
timestamp 1753449410
transform 1 0 10260 0 1 1032
box -446 -260 446 260
<< labels >>
flabel metal1 9386 938 9586 1138 0 FreeSans 256 0 0 0 Ibias
port 6 nsew default input
flabel metal1 9410 554 9610 754 0 FreeSans 256 0 0 0 VSS
port 3 nsew
flabel metal1 9378 3084 9578 3284 0 FreeSans 256 0 0 0 VDD
port 4 nsew
flabel metal1 10934 282 11134 482 0 FreeSans 256 0 0 0 V+
port 1 nsew
flabel metal1 10138 280 10338 480 0 FreeSans 256 0 0 0 V-
port 2 nsew default input
flabel metal1 11898 294 12098 494 0 FreeSans 256 0 0 0 Vout
port 5 nsew
<< end >>
