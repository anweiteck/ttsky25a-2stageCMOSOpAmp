* NGSPICE file created from 2stageCMOSOpAmp_parax.ext - technology: sky130A

.subckt 2stageCMOSOpAmp_parax V+ V- VSS VDD Vout Ibias
X0 VDD.t3 a_9954_2525# a_10740_2525# VDD.t2 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2.5
**devattr s=11600,516 d=11600,516
X1 VDD.t5 a_10740_2525# Vout.t1 VDD.t4 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0 ps=0 w=20 l=2.5
**devattr s=232000,8116 d=232000,8116
X2 a_10740_2525# Vout.t0 sky130_fd_pr__cap_mim_m3_1 l=20 w=20
X3 VSS.t6 Ibias.t2 Vout.t2 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=5 l=2.5
**devattr s=58000,2116 d=58000,2116
X4 a_10514_1672# V-.t0 a_9954_2525# VSS.t7 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.696 as=0.29 ps=2.58 w=1 l=2.5
**devattr s=11600,516 d=11600,516
X5 VDD.t1 a_9954_2525# a_9954_2525# VDD.t0 sky130_fd_pr__pfet_01v8 ad=0 pd=0 as=0.29 ps=2.58 w=1 l=2.5
**devattr s=11600,516 d=11600,516
X6 a_10514_1672# V+.t0 a_10740_2525# VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.696 as=0.29 ps=2.58 w=1 l=2.5
**devattr s=11600,516 d=11600,516
X7 VSS.t4 Ibias.t3 a_10514_1672# VSS.t3 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0.145 ps=1.348 w=0.5 l=2.5
**devattr s=5800,316 d=5800,316
X8 VSS.t2 Ibias.t0 Ibias.t1 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0 pd=0 as=0 ps=0 w=0.5 l=2.5
**devattr s=5800,316 d=5800,316
R0 VDD.n14 VDD.n12 8971.76
R1 VDD.n17 VDD.n11 8971.76
R2 VDD.n23 VDD.n8 2265.88
R3 VDD.n31 VDD.n4 2265.88
R4 VDD.n21 VDD.n3 1387.06
R5 VDD.n31 VDD.n3 1387.06
R6 VDD.n23 VDD.n6 1387.06
R7 VDD.n29 VDD.n6 1387.06
R8 VDD.n13 VDD.n9 956.989
R9 VDD.n13 VDD.n10 956.989
R10 VDD.n18 VDD.n10 956.989
R11 VDD.n25 VDD.n3 878.823
R12 VDD.n25 VDD.n6 878.823
R13 VDD.t2 VDD.n5 585.188
R14 VDD.t0 VDD.n5 585.188
R15 VDD.n19 VDD.n9 495.938
R16 VDD.n30 VDD.n4 480.914
R17 VDD.n22 VDD.n8 480.914
R18 VDD.n28 VDD.n2 241.695
R19 VDD.n24 VDD.n7 235.379
R20 VDD.n35 VDD.t1 233.118
R21 VDD.n0 VDD.t3 228.55
R22 VDD.n19 VDD.n18 151.861
R23 VDD.n27 VDD.n24 147.953
R24 VDD.n28 VDD.n27 147.953
R25 VDD.n32 VDD.n2 107.486
R26 VDD.n20 VDD.n19 106.236
R27 VDD.n26 VDD.n1 93.7417
R28 VDD.n27 VDD.n26 93.7417
R29 VDD.n16 VDD.n12 86.1255
R30 VDD.n15 VDD.n11 86.1255
R31 VDD.n19 VDD.n7 60.4449
R32 VDD.n8 VDD.n7 30.8338
R33 VDD.n4 VDD.n2 30.8338
R34 VDD.n26 VDD.n25 30.8338
R35 VDD.n25 VDD.n5 30.8338
R36 VDD.n14 VDD.n13 20.5561
R37 VDD.n18 VDD.n17 20.5561
R38 VDD.n29 VDD.n28 20.5561
R39 VDD.n24 VDD.n23 20.5561
R40 VDD.n23 VDD.t2 20.5561
R41 VDD.n21 VDD.n20 20.5561
R42 VDD.n32 VDD.n31 20.5561
R43 VDD.n31 VDD.t0 20.5561
R44 VDD.n17 VDD.n16 20.3127
R45 VDD.n15 VDD.n14 20.3127
R46 VDD.n30 VDD.n29 16.0482
R47 VDD.n22 VDD.n21 16.0482
R48 VDD.n0 VDD.t5 15.2715
R49 VDD.n20 VDD.n1 13.7448
R50 VDD.n33 VDD.n32 12.2759
R51 VDD.t2 VDD.n22 4.36374
R52 VDD.t0 VDD.n30 4.36374
R53 VDD.n11 VDD.n9 3.03329
R54 VDD.n12 VDD.n10 3.03329
R55 VDD.n33 VDD.n1 1.46935
R56 VDD VDD.n35 0.979373
R57 VDD.n34 VDD.n0 0.725365
R58 VDD.n34 VDD.n33 0.358192
R59 VDD.n16 VDD.t4 0.198323
R60 VDD.t4 VDD.n15 0.198323
R61 VDD.n35 VDD.n34 0.0577183
R62 Vout.n1 Vout.t2 17.3591
R63 Vout.n0 Vout.t1 12.4305
R64 Vout.n0 Vout.t0 5.96113
R65 Vout Vout.n1 2.08622
R66 Vout.n1 Vout.n0 1.82199
R67 Ibias.n5 Ibias.t1 229.112
R68 Ibias.n1 Ibias.t2 39.6502
R69 Ibias.n2 Ibias.t3 33.1654
R70 Ibias.t3 Ibias.n0 33.1654
R71 Ibias.n4 Ibias.t0 16.5847
R72 Ibias.n6 Ibias 2.08383
R73 Ibias.n1 Ibias.n0 1.059
R74 Ibias.n4 Ibias.n3 0.984715
R75 Ibias.n6 Ibias.n5 0.217566
R76 Ibias.n5 Ibias.n4 0.144319
R77 Ibias.n2 Ibias.n1 0.066125
R78 Ibias.n3 Ibias.n0 0.0412609
R79 Ibias.n3 Ibias.n2 0.00635938
R80 Ibias Ibias.n6 0.00274551
R81 VSS.n43 VSS.n42 353802
R82 VSS.n28 VSS.n25 5985.32
R83 VSS.n40 VSS.n24 5985.32
R84 VSS.n40 VSS.n25 5985.32
R85 VSS.n34 VSS.n32 3667.68
R86 VSS.n34 VSS.n33 3667.68
R87 VSS.n49 VSS.n12 3667.68
R88 VSS.n50 VSS.n12 3667.68
R89 VSS.n55 VSS.n3 3377.97
R90 VSS.n56 VSS.n3 3377.97
R91 VSS.n44 VSS.n19 3377.97
R92 VSS.n44 VSS.n20 3377.97
R93 VSS.n32 VSS.n16 2277.09
R94 VSS.n49 VSS.n16 2277.09
R95 VSS.n33 VSS.n11 2277.09
R96 VSS.n50 VSS.n11 2277.09
R97 VSS.n55 VSS.n6 2277.09
R98 VSS.n19 VSS.n6 2277.09
R99 VSS.n56 VSS.n4 2277.09
R100 VSS.n20 VSS.n4 2277.09
R101 VSS.n16 VSS.n15 1390.59
R102 VSS.n15 VSS.n11 1390.59
R103 VSS.n41 VSS.n23 1135.48
R104 VSS.n13 VSS.n6 1100.88
R105 VSS.n13 VSS.n4 1100.88
R106 VSS.n22 VSS.t0 836.559
R107 VSS.t3 VSS.n5 836.559
R108 VSS.t7 VSS.n14 836.559
R109 VSS.n21 VSS.t1 836.559
R110 VSS.n28 VSS.n27 759.684
R111 VSS.n42 VSS.n41 468.817
R112 VSS.n30 VSS.n29 388.906
R113 VSS.n42 VSS.t5 376.344
R114 VSS.n36 VSS.n30 368.565
R115 VSS.n29 VSS.n26 259.104
R116 VSS.n35 VSS.n31 238.306
R117 VSS.n0 VSS.t4 229.549
R118 VSS.n60 VSS.t2 229.538
R119 VSS.n48 VSS.n47 179.685
R120 VSS.n31 VSS.n17 147.953
R121 VSS.n48 VSS.n17 147.953
R122 VSS.n37 VSS.n3 146.25
R123 VSS.n22 VSS.n3 146.25
R124 VSS.n13 VSS.n9 146.25
R125 VSS.n14 VSS.n13 146.25
R126 VSS.n45 VSS.n44 146.25
R127 VSS.n44 VSS.n43 146.25
R128 VSS.n15 VSS.n8 117.001
R129 VSS.n15 VSS.n5 117.001
R130 VSS.n47 VSS.n12 117.001
R131 VSS.n21 VSS.n12 117.001
R132 VSS.n35 VSS.n34 117.001
R133 VSS.n34 VSS.n23 117.001
R134 VSS.n17 VSS.n8 90.3534
R135 VSS.n53 VSS.n8 90.3534
R136 VSS.n36 VSS.n35 90.3534
R137 VSS.n9 VSS.n2 71.5299
R138 VSS.n52 VSS.n9 70.777
R139 VSS.n32 VSS.n31 65.0005
R140 VSS.n32 VSS.t0 65.0005
R141 VSS.n49 VSS.n48 65.0005
R142 VSS.t7 VSS.n49 65.0005
R143 VSS.n26 VSS.n25 65.0005
R144 VSS.n25 VSS.t5 65.0005
R145 VSS.n30 VSS.n24 65.0005
R146 VSS.n55 VSS.n54 65.0005
R147 VSS.t3 VSS.n55 65.0005
R148 VSS.n19 VSS.n10 65.0005
R149 VSS.n19 VSS.t1 65.0005
R150 VSS.n51 VSS.n50 65.0005
R151 VSS.n50 VSS.t7 65.0005
R152 VSS.n33 VSS.n7 65.0005
R153 VSS.n33 VSS.t0 65.0005
R154 VSS.n20 VSS.n18 65.0005
R155 VSS.n20 VSS.t1 65.0005
R156 VSS.n57 VSS.n56 65.0005
R157 VSS.n56 VSS.t3 65.0005
R158 VSS.n27 VSS.n24 56.1412
R159 VSS.n29 VSS.n28 34.4123
R160 VSS.n40 VSS.n39 34.4123
R161 VSS.n41 VSS.n40 34.4123
R162 VSS.n45 VSS.n18 31.8499
R163 VSS.n46 VSS.n10 20.3492
R164 VSS.n0 VSS.t6 18.6429
R165 VSS.n57 VSS.n2 17.5893
R166 VSS.n18 VSS.n2 17.5893
R167 VSS.n26 VSS.n1 17.1124
R168 VSS.n54 VSS.n53 15.9595
R169 VSS.n52 VSS.n51 15.9595
R170 VSS.n38 VSS.n7 15.262
R171 VSS.n47 VSS.n46 12.191
R172 VSS.n58 VSS.n1 9.84665
R173 VSS.n46 VSS.n45 9.54971
R174 VSS.n23 VSS.n22 8.60265
R175 VSS.t3 VSS.t0 8.60265
R176 VSS.n14 VSS.n5 8.60265
R177 VSS.t7 VSS.t1 8.60265
R178 VSS.n43 VSS.n21 8.60265
R179 VSS.n27 VSS.t5 8.25109
R180 VSS.n38 VSS.n37 7.78001
R181 VSS.n37 VSS.n1 7.53124
R182 VSS.n58 VSS.n57 6.98232
R183 VSS.n39 VSS.n38 2.30721
R184 VSS.n39 VSS.n36 1.2217
R185 VSS VSS.n60 0.785005
R186 VSS.n60 VSS.n59 0.366479
R187 VSS.n54 VSS.n7 0.164603
R188 VSS.n53 VSS.n52 0.164603
R189 VSS.n51 VSS.n10 0.164603
R190 VSS.n59 VSS.n0 0.142897
R191 VSS.n59 VSS.n58 0.113915
R192 V- V-.t0 22.0581
R193 V+ V+.t0 22.0601
C0 Ibias a_9954_2525# 0.02164f
C1 V- a_10740_2525# 0.02337f
C2 Ibias a_10514_1672# 0.4269f
C3 a_10514_1672# a_9954_2525# 0.01029f
C4 Ibias VDD 0.03327f
C5 VDD a_9954_2525# 4.20596f
C6 VDD a_10514_1672# 0.03752f
C7 Ibias Vout 1.40938f
C8 Vout a_9954_2525# 0.07331f
C9 Ibias V+ 0.57534f
C10 a_9954_2525# V+ 0.06406f
C11 Vout a_10514_1672# 0.04417f
C12 Ibias a_10740_2525# 0.07752f
C13 a_10514_1672# V+ 0.77894f
C14 VDD Vout 2.92558f
C15 a_9954_2525# a_10740_2525# 0.64358f
C16 VDD V+ 0.02101f
C17 a_10514_1672# a_10740_2525# 0.23458f
C18 VDD a_10740_2525# 5.59104f
C19 Vout V+ 0.13377f
C20 Ibias V- 0.67f
C21 Vout a_10740_2525# 4.1443f
C22 V- a_9954_2525# 0.18797f
C23 V+ a_10740_2525# 0.14311f
C24 a_10514_1672# V- 0.2238f
C25 VDD V- 0.02203f
C26 Vout V- 0.00104f
C27 V- V+ 0.10701f
C28 Ibias VSS 8.48334f
C29 V+ VSS 2.32487f
C30 V- VSS 2.6456f
C31 Vout VSS 11.5548f
C32 VDD VSS 21.77651f
C33 a_10514_1672# VSS 1.16372f
C34 a_10740_2525# VSS 1.76783f
C35 a_9954_2525# VSS 1.75659f
C36 Vout.t1 VSS 0.09257f
C37 Vout.t0 VSS 6.30849f
C38 Vout.n0 VSS 0.29187f
C39 Vout.t2 VSS 0.01931f
C40 Vout.n1 VSS 0.22426f
C41 VDD.t3 VSS 0.0148f
C42 VDD.t5 VSS 0.68932f
C43 VDD.n0 VSS 1.90938f
C44 VDD.n1 VSS 0.1152f
C45 VDD.n2 VSS 0.0217f
C46 VDD.n3 VSS 0.02418f
C47 VDD.n4 VSS 0.23875f
C48 VDD.n5 VSS 0.34454f
C49 VDD.n6 VSS 0.02418f
C50 VDD.n7 VSS 0.02045f
C51 VDD.n8 VSS 0.23875f
C52 VDD.n9 VSS 0.09377f
C53 VDD.n10 VSS 0.11901f
C54 VDD.n11 VSS 1.58759f
C55 VDD.n12 VSS 1.58759f
C56 VDD.n13 VSS 0.1201f
C57 VDD.n14 VSS 0.1201f
C58 VDD.t4 VSS 2.50251f
C59 VDD.n17 VSS 0.1201f
C60 VDD.n18 VSS 0.0809f
C61 VDD.n19 VSS 0.70009f
C62 VDD.n20 VSS 0.28896f
C63 VDD.n21 VSS 0.02449f
C64 VDD.t2 VSS 0.35548f
C65 VDD.n23 VSS 0.02449f
C66 VDD.n24 VSS 0.02441f
C67 VDD.n25 VSS 0.01163f
C68 VDD.n26 VSS 0.01163f
C69 VDD.n27 VSS 0.02418f
C70 VDD.n28 VSS 0.02449f
C71 VDD.n29 VSS 0.02449f
C72 VDD.t0 VSS 0.35548f
C73 VDD.n31 VSS 0.02449f
C74 VDD.n32 VSS 0.18984f
C75 VDD.n33 VSS 0.09882f
C76 VDD.n34 VSS 0.08777f
C77 VDD.t1 VSS 0.01702f
C78 VDD.n35 VSS 0.30532f
.ends

